module dequan
#(
parameter IN_WIDTH = 12
)
(
input clk,
input Q_mode, // 0: Y, 1: U, V
input [2:0] read_addr,
input signed [IN_WIDTH-1:0] in0,
input signed [IN_WIDTH-1:0] in1,
input signed [IN_WIDTH-1:0] in2,
input signed [IN_WIDTH-1:0] in3,
input signed [IN_WIDTH-1:0] in4,
input signed [IN_WIDTH-1:0] in5,
input signed [IN_WIDTH-1:0] in6,
input signed [IN_WIDTH-1:0] in7,

//output reg [2:0] reg_waddr,
output [8*IN_WIDTH-1:0] out
);

//reg [2:0] reg_waddr_last;

reg signed [IN_WIDTH-1:0] i0, i1, i2, i3, i4, i5, i6, i7;

// quantized table
reg signed [8:0] QT0, QT1, QT2, QT3, QT4, QT5, QT6, QT7;
reg signed [8:0] QT00, QT11, QT22, QT33, QT44, QT55, QT66, QT77;
// quantized output
reg signed [IN_WIDTH+9-1:0] Q00, Q11, Q22, Q33, Q44, Q55, Q66, Q77;

assign out = {Q77[IN_WIDTH-1:0], Q66[IN_WIDTH-1:0], Q55[IN_WIDTH-1:0], Q44[IN_WIDTH-1:0], Q33[IN_WIDTH-1:0], Q22[IN_WIDTH-1:0],
              Q11[IN_WIDTH-1:0], Q00[IN_WIDTH-1:0]};


always @(posedge clk)
begin
  
//  reg_waddr_last <= read_addr;
//  reg_waddr <= reg_waddr_last;

  Q00        <= QT00 * i0;
  Q11        <= QT11 * i1;
  Q22        <= QT22 * i2;
  Q33        <= QT33 * i3;
  Q44        <= QT44 * i4;
  Q55        <= QT55 * i5;
  Q66        <= QT66 * i6;
  Q77        <= QT77 * i7;
  i0 <= in0;
  i1 <= in1;
  i2 <= in2;
  i3 <= in3;
  i4 <= in4;
  i5 <= in5;
  i6 <= in6;
  i7 <= in7;
  QT00 <= QT0;
  QT11 <= QT1;
  QT22 <= QT2;
  QT33 <= QT3;
  QT44 <= QT4;
  QT55 <= QT5;
  QT66 <= QT6;
  QT77 <= QT7;
end

always @*
begin
  case ({~Q_mode, read_addr}) // synopsys parallel_case
    4'b0000: begin
      QT0 = 9'd16;  // 1/16 = 0.062500 = 000010000 = 0.0625
      QT1 = 9'd11;  // 1/11 = 0.090909 = 000010111 = 0.08984375
      QT2 = 9'd10;  // 1/10 = 0.100000 = 000011010 = 0.1015625
      QT3 = 9'd16;  // 1/16 = 0.062500 = 000010000 = 0.0625
      QT4 = 9'd23;  // 1/24 = 0.041667 = 000001011 = 0.04296875
      QT5 = 9'd43;  // 1/40 = 0.025000 = 000000110 = 0.0234375
      QT6 = 9'd51;  // 1/51 = 0.019607 = 000000101 = 0.01953125
      QT7 = 9'd64;  // 1/61 = 0.016393 = 000000100 = 0.015625
    end
    4'b0001: begin
      QT0 = 9'd12;  // 1/12 = 0.083333 = 000010101 = 0.08203125
      QT1 = 9'd12;  // 1/12 = 0.083333 = 000010101 = 0.08203125
      QT2 = 9'd14;  // 1/14 = 0.071428 = 000010010 = 0.0703125
      QT3 = 9'd20;  // 1/19 = 0.052631 = 000001101 = 0.05078125
      QT4 = 9'd26;  // 1/26 = 0.038461 = 000001010 = 0.0390625
      QT5 = 9'd64;  // 1/58 = 0.017241 = 000000100 = 0.015625
      QT6 = 9'd64;  // 1/60 = 0.016667 = 000000100 = 0.015625
      QT7 = 9'd51;  // 1/55 = 0.018181 = 000000101 = 0.01953125
    end
    4'b0010: begin
      QT0 = 9'd14;  // 1/14 = 0.071428 = 000010010 = 0.0703125
      QT1 = 9'd13;  // 1/13 = 0.076923 = 000010100 = 0.078125
      QT2 = 9'd16;  // 1/16 = 0.062500 = 000010000 = 0.0625 
      QT3 = 9'd23;  // 1/24 = 0.041667 = 000001011 = 0.04296875
      QT4 = 9'd43;  // 1/40 = 0.025000 = 000000110 = 0.0234375
      QT5 = 9'd64;  // 1/57 = 0.017543 = 000000100 = 0.015625
      QT6 = 9'd64;  // 1/69 = 0.014492 = 000000100 = 0.015625
      QT7 = 9'd51;  // 1/56 = 0.017857 = 000000101 = 0.01953125
    end
    4'b0011: begin
      QT0 = 9'd14;  // 1/14 = 0.071428 = 000010010 = 0.0703125
      QT1 = 9'd17;  // 1/17 = 0.058823 = 000001111 = 0.05859375
      QT2 = 9'd21;  // 1/22 = 0.045454 = 000001100 = 0.046875
      QT3 = 9'd28;  // 1/29 = 0.034482 = 000001001 = 0.03515625
      QT4 = 9'd51;  // 1/51 = 0.019607 = 000000101 = 0.01953125
      QT5 = 9'd85;  // 1/87 = 0.011494 = 000000011 = 0.01171875
      QT6 = 9'd85;  // 1/80 = 0.012500 = 000000011 = 0.01171875
      QT7 = 9'd64;  // 1/62 = 0.016129 = 000000100 = 0.015625
    end
    4'b0100: begin
      QT0 = 9'd18;  // 1/18 = 0.055556 = 000001110 = 0.0546875
      QT1 = 9'd21;  // 1/22 = 0.045454 = 000001100 = 0.046875
      QT2 = 9'd37;  // 1/37 = 0.027027 = 000000111 = 0.02734375
      QT3 = 9'd51;  // 1/56 = 0.017857 = 000000101 = 0.01953125 
      QT4 = 9'd64;  // 1/68 = 0.014705 = 000000100 = 0.015625
      QT5 = 9'd128;  // 1/109 = 0.009174 = 000000010 = 0.0078125
      QT6 = 9'd128;  // 1/103 = 0.009708 = 000000010 = 0.0078125
      QT7 = 9'd85;  // 1/77 = 0.012987 = 000000011 = 0.01171875
    end
    4'b0101: begin
      QT0 = 9'd23;  // 1/24 = 0.041667 = 000001011 = 0.04296875
      QT1 = 9'd37;  // 1/35 = 0.028571 = 000000111 = 0.02734375
      QT2 = 9'd51;  // 1/55 = 0.018181 = 000000101 = 0.01953125
      QT3 = 9'd64;  // 1/64 = 0.015625 = 000000100 = 0.015625
      QT4 = 9'd85;  // 1/81 = 0.012345 = 000000011 = 0.01171875
      QT5 = 9'd128;  // 1/104 = 0.009615 = 000000010 = 0.0078125
      QT6 = 9'd128;  // 1/113 = 0.008849 = 000000010 = 0.0078125
      QT7 = 9'd85;  // 1/92 = 0.010869 = 000000011 = 0.01171875
    end
    4'b0110: begin
      QT0 = 9'd51;  // 1/49 = 0.020408 = 000000101 = 0.01953125
      QT1 = 9'd64;  // 1/64 = 0.015625 = 000000100 = 0.015625
      QT2 = 9'd85;  // 1/78 = 0.012820 = 000000011 = 0.01171875
      QT3 = 9'd85;  // 1/87 = 0.011494 = 000000011 = 0.01171875
      QT4 = 9'd128;  // 1/103 = 0.009708 = 000000010 = 0.0078125
      QT5 = 9'd128;  // 1/121 = 0.008264 = 000000010 = 0.0078125 
      QT6 = 9'd128;  // 1/120 = 0.008333 = 000000010 = 0.0078125
      QT7 = 9'd85;  // 1/101 = 0.009901 = 000000011 = 0.01171875
    end
    4'b0111: begin
      QT0 = 9'd64;  // 1/72 = 0.013888 = 000000100 = 0.015625
      QT1 = 9'd85;  // 1/92 = 0.010869 = 000000011 = 0.01171875
      QT2 = 9'd85;  // 1/95 = 0.010526 = 000000011 = 0.01171875
      QT3 = 9'd85;  // 1/98 = 0.010204 = 000000011 = 0.01171875
      QT4 = 9'd128;  // 1/112 = 0.008928 = = 000000010 = 0.0078125
      QT5 = 9'd85;  // 1/100 = 0.010000 = 000000011 = 0.01171875
      QT6 = 9'd128;  // 1/103 = 0.009708 = 000000010 = 0.0078125
      QT7 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
    end
    4'b1000: begin
      QT0 = 9'd17;  // 1/17 = 0.058823 = 000001111 = 0.05859375
      QT1 = 9'd18;  // 1/18 = 0.055556 = 000001110 = 0.0546875
      QT2 = 9'd23;  // 1/24 = 0.041667 = 000001011 = 0.04296875
      QT3 = 9'd51;  // 1/47 = 0.021276 = 000000101 = 0.01953125
      QT4 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT5 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT6 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT7 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
    end
    4'b1001: begin
      QT0 = 9'd18;  // 1/18 = 0.055556 = 000001110 = 0.0546875
      QT1 = 9'd21;  // 1/21 = 0.047619 = 000001100 = 0.046875
      QT2 = 9'd26;  // 1/26 = 0.038461 = 000001010 = 0.0390625
      QT3 = 9'd64;  // 1/66 = 0.015152 = 000000100 = 0.015625
      QT4 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT5 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT6 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT7 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
    end
    4'b1010: begin
      QT0 = 9'd23;  // 1/24 = 0.041667 = 000001011 = 0.04296875
      QT1 = 9'd26;  // 1/26 = 0.038461 = 000001010 = 0.0390625
      QT2 = 9'd51;  // 1/56 = 0.017857 = 000000101 = 0.01953125
      QT3 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT4 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT5 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT6 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT7 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
    end
    4'b1011: begin
      QT0 = 9'd51;  // 1/47 = 0.021276 = 000000101 = 0.01953125
      QT1 = 9'd64;  // 1/66 = 0.015152 = 000000100 = 0.015625
      QT2 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT3 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT4 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT5 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT6 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT7 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
    end
    4'b1100: begin
      QT0 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT1 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT2 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT3 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT4 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT5 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT6 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT7 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
    end
    4'b1101: begin
      QT0 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT1 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT2 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT3 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT4 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT5 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT6 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT7 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
    end
    4'b1110: begin
      QT0 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT1 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT2 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT3 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT4 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT5 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT6 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT7 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
    end
    4'b1111: begin
      QT0 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT1 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT2 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT3 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT4 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875 
      QT5 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT6 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
      QT7 = 9'd85;  // 1/99 = 0.010101 = 000000011 = 0.01171875
    end
    default: begin
      QT0 = 9'd0;
      QT1 = 9'd0; 
      QT2 = 9'd0;
      QT3 = 9'd0;
      QT4 = 9'd0; 
      QT5 = 9'd0; 
      QT6 = 9'd0; 
      QT7 = 9'd0;
    end
  endcase
end


endmodule
